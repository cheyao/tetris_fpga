module position_counter (
    input [9:0] sq2, sq0,
    output reg [4:0] pos1, pos0
);
    wire [19:0] act_row;

	generate
    genvar i;
	for(i = 0; i<20; i = i+1) begin : bc
		assign act_row[i] = sq0 <= 10'd60 + 20 * i ;
	end
	endgenerate

	always @* begin

        case(sq2)
		10'd240: pos0 = 5'd0;
		10'd260: pos0 = 5'd1;
		10'd280: pos0 = 5'd2;
		10'd300: pos0 = 5'd3;
		10'd320: pos0 = 5'd4;
		10'd340: pos0 = 5'd5;
		10'd360: pos0 = 5'd6;
		10'd380: pos0 = 5'd7;
		10'd400: pos0 = 5'd8;
		10'd420: pos0 = 5'd9;
		default: pos0 = 5'd10;
	    endcase

        casez(act_row)
		20'b???????????????????1: pos1 = 5'd0;
		20'b??????????????????10: pos1 = 5'd1;
		20'b?????????????????100: pos1 = 5'd2;
		20'b????????????????1000: pos1 = 5'd3;
		20'b???????????????10000: pos1 = 5'd4;
		20'b??????????????100000: pos1 = 5'd5;
		20'b?????????????1000000: pos1 = 5'd6;
		20'b????????????10000000: pos1 = 5'd7;
		20'b???????????100000000: pos1 = 5'd8;
		20'b??????????1000000000: pos1 = 5'd9;
		20'b?????????10000000000: pos1 = 5'd10;
		20'b????????100000000000: pos1 = 5'd11;
		20'b???????1000000000000: pos1 = 5'd12;
		20'b??????10000000000000: pos1 = 5'd13;
		20'b?????100000000000000: pos1 = 5'd14;
		20'b????1000000000000000: pos1 = 5'd15;
		20'b???10000000000000000: pos1 = 5'd16;
		20'b??100000000000000000: pos1 = 5'd17;
		20'b?1000000000000000000: pos1 = 5'd18;
		20'b10000000000000000000: pos1 = 5'd19;
		default: pos1 = 5'd0;
	    endcase
    end
endmodule