// clock_divider.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module clock_divider (
		output wire  clk_clk,        //      clk.clk
		input  wire  clk_in_clk,     //   clk_in.clk
		input  wire  reset_in_reset  // reset_in.reset
	);

	clock_divider_pll_0 pll_0 (
		.refclk   (clk_in_clk),     //  refclk.clk
		.rst      (reset_in_reset), //   reset.reset
		.outclk_0 (clk_clk),        // outclk0.clk
		.locked   ()                // (terminated)
	);

endmodule
